`ifndef src__slash__snow64_alu_defines_header_sv
`define src__slash__snow64_alu_defines_header_sv

// src/snow64_alu_defines.header.sv

`include "src/misc_defines.header.sv"

`define WIDTH__SNOW64_ALU_OPER 4
`define MSB_POS__SNOW64_ALU_OPER `WIDTH2MP(`WIDTH__SNOW64_ALU_OPER)

`define WIDTH__SNOW64_ALU_TYPE_SIZE 2
`define MSB_POS__SNOW64_ALU_TYPE_SIZE \
	`WIDTH2MP(`WIDTH__SNOW64_ALU_TYPE_SIZE)

`define WIDTH__SNOW64_ALU_BREAK_INDEX 2
`define MSB_POS__SNOW64_ALU_BREAK_INDEX \
	`WIDTH2MP(`WIDTH__SNOW64_ALU_BREAK_INDEX)

`define WIDTH__SNOW64_ALU_64_DATA_INOUT 64
`define MSB_POS__SNOW64_ALU_64_DATA_INOUT \
	`WIDTH2MP(`WIDTH__SNOW64_ALU_64_DATA_INOUT)
`define WIDTH__SNOW64_ALU_32_DATA_INOUT 32
`define MSB_POS__SNOW64_ALU_32_DATA_INOUT \
	`WIDTH2MP(`WIDTH__SNOW64_ALU_32_DATA_INOUT)
`define WIDTH__SNOW64_ALU_16_DATA_INOUT 16
`define MSB_POS__SNOW64_ALU_16_DATA_INOUT \
	`WIDTH2MP(`WIDTH__SNOW64_ALU_16_DATA_INOUT)
`define WIDTH__SNOW64_ALU_8_DATA_INOUT 8
`define MSB_POS__SNOW64_ALU_8_DATA_INOUT \
	`WIDTH2MP(`WIDTH__SNOW64_ALU_8_DATA_INOUT)

`define WIDTH__SNOW64_SUB_ALU_DATA_INOUT 8
`define MSB_POS__SNOW64_SUB_ALU_DATA_INOUT \
	`WIDTH2MP(`WIDTH__SNOW64_SUB_ALU_DATA_INOUT)

`define WIDTH__SNOW64_SUB_ALU_INDEX $clog2(64 / 8)
`define MSB_POS__SNOW64_SUB_ALU_INDEX \
	`WIDTH2MP(`WIDTH__SNOW64_SUB_ALU_INDEX)

`define WIDTH__SNOW64_ALU_NUM_8_BIT_SUB_ALUS $clog2(64 / 8)
`define MSB_POS__SNOW64_ALU_NUM_8_BIT_SUB_ALUS \
	`WIDTH2MP(`WIDTH__SNOW64_ALU_NUM_8_BIT_SUB_ALUS)

`define WIDTH__SNOW64_ALU_NUM_16_BIT_SUB_ALUS $clog2(64 / 16)
`define MSB_POS__SNOW64_ALU_NUM_16_BIT_SUB_ALUS \
	`WIDTH2MP(`WIDTH__SNOW64_ALU_NUM_16_BIT_SUB_ALUS)

`define WIDTH__SNOW64_ALU_NUM_32_BIT_SUB_ALUS $clog2(64 / 32)
`define MSB_POS__SNOW64_ALU_NUM_32_BIT_SUB_ALUS \
	`WIDTH2MP(`WIDTH__SNOW64_ALU_NUM_32_BIT_SUB_ALUS)

`endif		// src__slash__snow64_alu_defines_header_sv
