`ifndef src__slash__snow64_memory_access_via_fifos_defines_header_sv
`define src__slash__snow64_memory_access_via_fifos_defines_header_sv

// src/snow64_memory_access_via_fifos_defines.header.sv

//`include "src/misc_defines.header.sv"
`include "src/snow64_cpu_defines.header.sv"
`include "src/snow64_lar_file_defines.header.sv"



`endif		// src__slash__snow64_memory_access_via_fifos_defines_header_sv
