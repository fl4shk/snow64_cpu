`ifndef src__slash__snow64_alu_defines_header_sv
`define src__slash__snow64_alu_defines_header_sv

// src/snow64_alu_defines.header.sv

`include "src/misc_defines.header.sv"

`define WIDTH__SNOW64_ALU_OPER 4
`define MSB_POS__SNOW64_ALU_OPER `WIDTH2MP(`WIDTH__SNOW64_ALU_OPER)

`define WIDTH__SNOW64_SUB_ALU_OUT_SLT_8 8
`define MSB_POS__SNOW64_SUB_ALU_OUT_SLT_8 \
	`WIDTH2MP(`WIDTH__SNOW64_SUB_ALU_OUT_SLT_8)
`define WIDTH__SNOW64_SUB_ALU_OUT_SLT_16 4
`define MSB_POS__SNOW64_SUB_ALU_OUT_SLT_16 \
	`WIDTH2MP(`WIDTH__SNOW64_SUB_ALU_OUT_SLT_16)
`define WIDTH__SNOW64_SUB_ALU_OUT_SLT_32 2
`define MSB_POS__SNOW64_SUB_ALU_OUT_SLT_32 \
	`WIDTH2MP(`WIDTH__SNOW64_SUB_ALU_OUT_SLT_32)
`define WIDTH__SNOW64_SUB_ALU_OUT_SLT_64 1
`define MSB_POS__SNOW64_SUB_ALU_OUT_SLT_64 \
	`WIDTH2MP(`WIDTH__SNOW64_SUB_ALU_OUT_SLT_64)



`define WIDTH__SNOW64_SUB_ALU_DATA_INOUT 8
`define MSB_POS__SNOW64_SUB_ALU_DATA_INOUT \
	`WIDTH2MP(`WIDTH__SNOW64_SUB_ALU_DATA_INOUT)

`define WIDTH__SNOW64_SUB_ALU_INDEX $clog2(64 / 8)
`define MSB_POS__SNOW64_SUB_ALU_INDEX \
	`WIDTH2MP(`WIDTH__SNOW64_SUB_ALU_INDEX)
//`define WIDTH__SNOW64_SUB_ALU_DATA_INOUT 16
//`define MSB_POS__SNOW64_SUB_ALU_DATA_INOUT \
//	`WIDTH2MP(`WIDTH__SNOW64_SUB_ALU_DATA_INOUT)
//
//`define WIDTH__SNOW64_SUB_ALU_INDEX $clog2(64 / 16)
//`define MSB_POS__SNOW64_SUB_ALU_INDEX \
//	`WIDTH2MP(`WIDTH__SNOW64_SUB_ALU_INDEX)

`define ARR_SIZE__SNOW64_ALU_SLICE_AND_EXTEND_OUT_DATA 8
`define LAST_INDEX__SNOW64_ALU_SLICE_AND_EXTEND_OUT_DATA \
	`ARR_SIZE_TO_LAST_INDEX(`ARR_SIZE__SNOW64_ALU_SLICE_AND_EXTEND_OUT_DATA)

`endif		// src__slash__snow64_alu_defines_header_sv
