`ifndef src__slash__snow64_operand_manager_defines_header_sv
`define src__slash__snow64_operand_manager_defines_header_sv

// src/snow64_operand_manager_defines.header.sv

`include "src/snow64_cpu_defines.header.sv"
`include "src/snow64_lar_file_defines.header.sv"

`endif		// src__slash__snow64_operand_manager_defines_header_sv
