`include "src/snow64_bfloat16_defines.header.sv"

//module Snow64BFloat16Add(input logic clk,
//	input PkgSnow64BFloat16::PortIn_Add in,
//	output PkgSnow64BFloat16::PortOut_Add out);
//
//endmodule
