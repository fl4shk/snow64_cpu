`ifndef src__slash__snow64_instr_cache_defines_header_sv
`define src__slash__snow64_instr_cache_defines_header_sv

// src/snow64_instr_cache_defines.header.sv

`include "src/misc_defines.header.sv"
`include "src/snow64_lar_file_defines.header.sv"
`include "src/snow64_instr_decoder_defines.header.sv"



// A single icache line is as long as a single LAR.
// This is done for simplicity purposes.
`define WIDTH__SNOW64_ICACHE_LINE_DATA `WIDTH__SNOW64_LAR_FILE_DATA
`define MSB_POS__SNOW64_ICACHE_LINE_DATA \
	`WIDTH2MP(`WIDTH__SNOW64_ICACHE_LINE_DATA)

`define WIDTH__SNOW64_ICACHE_LINE_PACKED_OUTER_DIM `WIDTH__SNOW64_INSTR
//`define WIDTH__SNOW64_ICACHE_LINE_PACKED_OUTER_DIM 64
//`define WIDTH__SNOW64_ICACHE_LINE_PACKED_OUTER_DIM 16
`define MSB_POS__SNOW64_ICACHE_LINE_PACKED_OUTER_DIM \
	`WIDTH2MP(`WIDTH__SNOW64_ICACHE_LINE_PACKED_OUTER_DIM)

`define WIDTH__SNOW64_ICACHE_LINE_PACKED_INNER_DIM \
	(`WIDTH__SNOW64_ICACHE_LINE_DATA \
	/ `WIDTH__SNOW64_ICACHE_LINE_PACKED_OUTER_DIM)
`define MSB_POS__SNOW64_ICACHE_LINE_PACKED_INNER_DIM \
	`WIDTH2MP(`WIDTH__SNOW64_ICACHE_LINE_PACKED_INNER_DIM)


// Max possible number of addresses whose data is stored.
`define WIDTH__SNOW64_ICACHE_EFFECTIVE_ADDR__BYTE_BASE_ADDR 15
`define MSB_POS__SNOW64_ICACHE_EFFECTIVE_ADDR__BYTE_BASE_ADDR \
	`WIDTH2MP(`WIDTH__SNOW64_ICACHE_EFFECTIVE_ADDR__BYTE_BASE_ADDR)




// An index into the line of data (select an instruction from the line of
// data)
`define WIDTH__SNOW64_ICACHE_EFFECTIVE_ADDR__LINE_INDEX \
	($clog2(`WIDTH__SNOW64_ICACHE_LINE_PACKED_INNER_DIM))
`define MSB_POS__SNOW64_ICACHE_EFFECTIVE_ADDR__LINE_INDEX \
	`WIDTH2MP(`WIDTH__SNOW64_ICACHE_EFFECTIVE_ADDR__LINE_INDEX)


`define WIDTH__SNOW64_ICACHE_LINE_BYTE_INDEX \
	$clog2(`WIDTH__SNOW64_ICACHE_LINE_PACKED_INNER_DIM)
`define MSB_POS__SNOW64_ICACHE_LINE_BYTE_INDEX \
	`WIDTH2MP(`WIDTH__SNOW64_ICACHE_LINE_BYTE_INDEX)

// Forcefully align addresses to width of instructions
// if outer index width is 8, WIDTH...DONT_CARE == 0
// if outer index width is 16, WIDTH...DONT_CARE == 1
// if outer index width is 32, WIDTH...DONT_CARE == 2
`define WIDTH__SNOW64_ICACHE_EFFECTIVE_ADDR__DONT_CARE \
	$clog2(`WIDTH__SNOW64_ICACHE_LINE_PACKED_OUTER_DIM / 8)
`define MSB_POS__SNOW64_ICACHE_EFFECTIVE_ADDR__DONT_CARE \
	`WIDTH2MP(`WIDTH__SNOW64_ICACHE_EFFECTIVE_ADDR__DONT_CARE)

// 32 kiB instruction cache
`define ARR_SIZE__SNOW64_ICACHE_NUM_LINES \
	((1 << `WIDTH__SNOW64_ICACHE_EFFECTIVE_ADDR__BYTE_BASE_ADDR) \
	/ (`WIDTH__SNOW64_ICACHE_LINE_DATA / 8))
`define LAST_INDEX__SNOW64_ICACHE_NUM_LINES \
	`ARR_SIZE_TO_LAST_INDEX(ARR_SIZE__SNOW64_ICACHE_NUM_LINES)

`define WIDTH__SNOW64_ICACHE_EFFECTIVE_ADDR__ARR_INDEX \
	$clog2(`ARR_SIZE__SNOW64_ICACHE_NUM_LINES)
`define MSB_POS__SNOW64_ICACHE_EFFECTIVE_ADDR__ARR_INDEX \
	`WIDTH2MP(`WIDTH__SNOW64_ICACHE_EFFECTIVE_ADDR__ARR_INDEX)

`define WIDTH__SNOW64_ICACHE_EFFECTIVE_ADDR__TAG \
	(`WIDTH__SNOW64_CPU_ADDR \
	- `WIDTH__SNOW64_ICACHE_EFFECTIVE_ADDR__ARR_INDEX \
	- `WIDTH__SNOW64_ICACHE_EFFECTIVE_ADDR__LINE_INDEX \
	- `WIDTH__SNOW64_ICACHE_EFFECTIVE_ADDR__DONT_CARE)
`define MSB_POS__SNOW64_ICACHE_EFFECTIVE_ADDR__TAG \
	`WIDTH2MP(`WIDTH__SNOW64_ICACHE_EFFECTIVE_ADDR__TAG)


`endif		// src__slash__snow64_instr_cache_defines_header_sv
