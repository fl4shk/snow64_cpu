`ifndef src__slash__snow64_alu_defines_header_sv
`define src__slash__snow64_alu_defines_header_sv

// src/snow64_alu_defines.header.sv

`include "src/misc_defines.header.sv"

`define WIDTH__SNOW64_CPU_ALU_OPER 4
`define MSB_POS__SNOW64_CPU_ALU_OPER `WIDTH2MP(`WIDTH__SNOW64_CPU_ALU_OPER)


`define WIDTH__SNOW64_CPU_ALU_64_DATA_INOUT 64
`define MSB_POS__SNOW64_CPU_ALU_64_DATA_INOUT \
	`WIDTH2MP(`WIDTH__SNOW64_CPU_ALU_64_DATA_INOUT)
`define WIDTH__SNOW64_CPU_ALU_32_DATA_INOUT 32
`define MSB_POS__SNOW64_CPU_ALU_32_DATA_INOUT \
	`WIDTH2MP(`WIDTH__SNOW64_CPU_ALU_32_DATA_INOUT)
`define WIDTH__SNOW64_CPU_ALU_16_DATA_INOUT 16
`define MSB_POS__SNOW64_CPU_ALU_16_DATA_INOUT \
	`WIDTH2MP(`WIDTH__SNOW64_CPU_ALU_16_DATA_INOUT)
`define WIDTH__SNOW64_CPU_ALU_8_DATA_INOUT 8
`define MSB_POS__SNOW64_CPU_ALU_8_DATA_INOUT \
	`WIDTH2MP(`WIDTH__SNOW64_CPU_ALU_8_DATA_INOUT)

`define WIDTH__SNOW64_CPU_ALU_SHIFT_DATA_INOUT 64
`define MSB_POS__SNOW64_CPU_ALU_SHIFT_DATA_INOUT \
	`WIDTH2MP(`WIDTH__SNOW64_CPU_ALU_SHIFT_DATA_INOUT)
`define WIDTH__SNOW64_CPU_ALU_SHIFT_AMOUNT 6
`define MSB_POS__SNOW64_CPU_ALU_SHIFT_AMOUNT \
	`WIDTH2MP(`WIDTH__SNOW64_CPU_ALU_SHIFT_AMOUNT)

`endif		// src__slash__snow64_alu_defines_header_sv
